library ieee;
use ieee.std_logic_1164.all;

package top_config is

  constant N : positive := 8;
  constant ADDR_WIDTH : integer := 8;

end package top_config;